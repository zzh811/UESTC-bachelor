module adjust_test(clk,reset,press,updwnout);
	
	input clk,reset,press;
	output updwnout;

	reg updwnout;
	reg [31:0]cnt;
	
//-----------------------------


//-----------------------------

endmodule
